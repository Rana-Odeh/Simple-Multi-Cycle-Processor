module instruction_memory(clk,addr,out);
    input [31:0] addr;
    output reg [31:0] out;
    reg [31:0] mem [0:1023];
	input clk;
    always @( posedge clk or addr) begin
       out = mem[addr];
    end	 
	 initial begin
        // Set instructions directly in the memory array
        mem[0] = 32'b00000000000001001000000000000000; //AND
        mem[1] = 32'b00000100000001001000000000000000; // ADD 
        mem[2] = 32'b00001000000001001000000000000000 ;	 // sub
		mem[3] = 32'b00001100000001000000000000000100; //andi
		mem[4] = 32'b00010000000001000000000000000100; //addi
		mem[5] = 32'b00010100000001000000000000000100 ;// lw 	
		mem[6] = 32'b00011000000001000000000000000100;// lw _poi  
		mem[7] = 32'b 00011100000001000000000000000100;// sw 
		mem[8] = 32'b00100000000001000000000000000100 ;// bgt  
		mem[9] = 32'b 00100100000001000000000000001100; // blt
		mem[10] = 32'b 00101000000001000000000000000100; // beq
		mem[11] = 32'b 00101100000001000000000000000100; // bne
		mem[12] = 32'b 00110000000000000000000000000100	; // jmp
		mem[13] = 32'b 00110100000000000000000000000100; // call  
		mem[14] = 32'b 00111000000000000000000000000000; //ret	  
		mem[15] = 32'b 00111100010000000000000000000000	; //push
		mem[16] = 32'b 01000000010000000000000000000000 ; // pop 
		
		
    end
endmodule